module Pong (
    input clk,
    input rst,
    inout wire PS2_DATA,
	inout wire PS2_CLK,
    output reg [63:0] layer1,
    output reg [63:0] layer2,
    output reg [63:0] layer3,
    output reg [63:0] layer4,
    output reg [63:0] layer5,
    output reg [63:0] layer6,
    output reg [63:0] layer7,
    output reg [63:0] layer8
);
    reg cube[7:0][7:0][7:0]; // x y z

    reg [2:0] A_pos_x = 3'd4;
    reg [2:0] A_pos_z = 3'd4;
    reg [2:0] next_A_pos_x;
    reg [2:0] next_A_pos_z;

    reg [2:0] B_pos_x = 3'd4;
    reg [2:0] B_pos_z = 3'd4;
    reg [2:0] next_B_pos_x;
    reg [2:0] next_B_pos_z;

    reg [2:0] ball_pos_x;
    reg [2:0] next_ball_pos_x;
    reg [2:0] prev_ball_pos_x;
    reg [2:0] ball_pos_y;
    reg [2:0] next_ball_pos_y;
    reg [2:0] prev_ball_pos_y;
    reg [2:0] ball_pos_z;
    reg [2:0] next_ball_pos_z;
    reg [2:0] prev_ball_pos_z;
    reg [2:0] delta_x;
    reg [2:0] next_delta_x;
    reg [2:0] delta_y;
    reg [2:0] next_delta_y;
    reg [2:0] delta_z;
    reg [2:0] next_delta_z;

    reg [3:0] A_score;
    reg [3:0] next_A_score;
    reg [3:0] B_score;
    reg [3:0] next_B_score;

    reg Pause;
    reg Next_Pause;

	wire [511:0] key_down;
	wire [8:0] last_change;
	wire been_ready;
    wire clk_div;
    wire clk_div_25;
    wire clk_div_26;

    reg [1:0] state;
    reg [1:0] Next_state;

    parameter ShowScore_1 = 2'b0;
    parameter ShowScore_2 = 2'b01;
    parameter Play = 2'b10;

    parameter A_Up      = 9'b0_0001_1101; // W => 1D
    parameter A_Down    = 9'b0_0001_1011; // S => 1B
    parameter A_Right   = 9'b0_0001_1100; // A => 1C
    parameter A_Left    = 9'b0_0010_0011; // D => 23
    parameter B_Up      = 9'b0_0111_0011; // 5 => 73
    parameter B_Down    = 9'b0_0111_0010; // 2 => 72
    parameter B_Left    = 9'b0_0110_1001; // 1 => 69
    parameter B_Right   = 9'b0_0111_1010; // 3 => 7A
    parameter Space     = 9'b0_0010_1001; // space => 29

    parameter pos = 1;
    parameter neg = -1;

	KeyboardDecoder key_de (
		.key_down(key_down),
		.last_change(last_change),
		.key_valid(been_ready),
		.PS2_DATA(PS2_DATA),
		.PS2_CLK(PS2_CLK),
		.rst(rst),
		.clk(clk)
	);

    clockDivider #(.n(25)) Clk26(clk, clk_div_26);
    clockDivider #(.n(24)) Clk25(clk, clk_div_25);

    assign clk_div = (A_score > 7 || B_score > 7)? clk_div_25 : clk_div_26;

    always @(posedge clk_div, posedge rst) begin
        if (rst) begin
            ball_pos_x <= 3'd4;
            ball_pos_y <= 3'd1;
            ball_pos_z <= 3'd4;
            delta_x <= 0;
            delta_y <= 1;
            delta_z <= 0;
            prev_ball_pos_x <= 3'd4;
            prev_ball_pos_y <= 3'd4;
            prev_ball_pos_z <= 3'd4;
            A_score <= 4'b0;
            B_score <= 4'b0;
            state <= Play;
        end
        else begin
            if (!Pause) begin
                prev_ball_pos_x <= ball_pos_x;
                prev_ball_pos_y <= ball_pos_y;
                prev_ball_pos_z <= ball_pos_z;
                ball_pos_x <= next_ball_pos_x;
                ball_pos_y <= next_ball_pos_y;
                ball_pos_z <= next_ball_pos_z;
                A_score <= next_A_score;
                B_score <= next_B_score;
                delta_x <= next_delta_x;
                delta_y <= next_delta_y;
                delta_z <= next_delta_z;
                state <= Next_state;
            end
        end
        
    end

    always @ (posedge clk, posedge rst) begin
		if (rst) begin
            A_pos_x <= 3'd4;
            A_pos_z <= 3'd4;
            B_pos_x <= 3'd4;
            B_pos_z <= 3'd4;
            layer1 <= 64'b0;
            layer2 <= 64'b0;
            layer3 <= 64'b0;
            layer4 <= 64'b0;
            layer5 <= 64'b0;
            layer6 <= 64'b0;
            layer7 <= 64'b0;
            layer8 <= 64'b0;
            Pause <= 1'b1;
            cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
            cube[0][1][0] <= 1'b0; cube[1][1][0] <= 1'b0; cube[2][1][0] <= 1'b0; cube[3][1][0] <= 1'b0; cube[4][1][0] <= 1'b0; cube[5][1][0] <= 1'b0; cube[6][1][0] <= 1'b0; cube[7][1][0] <= 1'b0; 
            cube[0][2][0] <= 1'b0; cube[1][2][0] <= 1'b0; cube[2][2][0] <= 1'b0; cube[3][2][0] <= 1'b0; cube[4][2][0] <= 1'b0; cube[5][2][0] <= 1'b0; cube[6][2][0] <= 1'b0; cube[7][2][0] <= 1'b0; 
            cube[0][3][0] <= 1'b0; cube[1][3][0] <= 1'b0; cube[2][3][0] <= 1'b0; cube[3][3][0] <= 1'b0; cube[4][3][0] <= 1'b0; cube[5][3][0] <= 1'b0; cube[6][3][0] <= 1'b0; cube[7][3][0] <= 1'b0;
            cube[0][4][0] <= 1'b0; cube[1][4][0] <= 1'b0; cube[2][4][0] <= 1'b0; cube[3][4][0] <= 1'b0; cube[4][4][0] <= 1'b0; cube[5][4][0] <= 1'b0; cube[6][4][0] <= 1'b0; cube[7][4][0] <= 1'b0; 
            cube[0][5][0] <= 1'b0; cube[1][5][0] <= 1'b0; cube[2][5][0] <= 1'b0; cube[3][5][0] <= 1'b0; cube[4][5][0] <= 1'b0; cube[5][5][0] <= 1'b0; cube[6][5][0] <= 1'b0; cube[7][5][0] <= 1'b0; 
            cube[0][6][0] <= 1'b0; cube[1][6][0] <= 1'b0; cube[2][6][0] <= 1'b0; cube[3][6][0] <= 1'b0; cube[4][6][0] <= 1'b0; cube[5][6][0] <= 1'b0; cube[6][6][0] <= 1'b0; cube[7][6][0] <= 1'b0;
            cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
            cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b0; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b0; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0; 
            cube[0][1][1] <= 1'b0; cube[1][1][1] <= 1'b0; cube[2][1][1] <= 1'b0; cube[3][1][1] <= 1'b0; cube[4][1][1] <= 1'b0; cube[5][1][1] <= 1'b0; cube[6][1][1] <= 1'b0; cube[7][1][1] <= 1'b0;
            cube[0][2][1] <= 1'b0; cube[1][2][1] <= 1'b0; cube[2][2][1] <= 1'b0; cube[3][2][1] <= 1'b0; cube[4][2][1] <= 1'b0; cube[5][2][1] <= 1'b0; cube[6][2][1] <= 1'b0; cube[7][2][1] <= 1'b0; 
            cube[0][3][1] <= 1'b0; cube[1][3][1] <= 1'b0; cube[2][3][1] <= 1'b0; cube[3][3][1] <= 1'b0; cube[4][3][1] <= 1'b0; cube[5][3][1] <= 1'b0; cube[6][3][1] <= 1'b0; cube[7][3][1] <= 1'b0; 
            cube[0][4][1] <= 1'b0; cube[1][4][1] <= 1'b0; cube[2][4][1] <= 1'b0; cube[3][4][1] <= 1'b0; cube[4][4][1] <= 1'b0; cube[5][4][1] <= 1'b0; cube[6][4][1] <= 1'b0; cube[7][4][1] <= 1'b0;
            cube[0][5][1] <= 1'b0; cube[1][5][1] <= 1'b0; cube[2][5][1] <= 1'b0; cube[3][5][1] <= 1'b0; cube[4][5][1] <= 1'b0; cube[5][5][1] <= 1'b0; cube[6][5][1] <= 1'b0; cube[7][5][1] <= 1'b0; 
            cube[0][6][1] <= 1'b0; cube[1][6][1] <= 1'b0; cube[2][6][1] <= 1'b0; cube[3][6][1] <= 1'b0; cube[4][6][1] <= 1'b0; cube[5][6][1] <= 1'b0; cube[6][6][1] <= 1'b0; cube[7][6][1] <= 1'b0; 
            cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b0; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0; 
            cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
            cube[0][1][2] <= 1'b0; cube[1][1][2] <= 1'b0; cube[2][1][2] <= 1'b0; cube[3][1][2] <= 1'b0; cube[4][1][2] <= 1'b0; cube[5][1][2] <= 1'b0; cube[6][1][2] <= 1'b0; cube[7][1][2] <= 1'b0; 
            cube[0][2][2] <= 1'b0; cube[1][2][2] <= 1'b0; cube[2][2][2] <= 1'b0; cube[3][2][2] <= 1'b0; cube[4][2][2] <= 1'b0; cube[5][2][2] <= 1'b0; cube[6][2][2] <= 1'b0; cube[7][2][2] <= 1'b0; 
            cube[0][3][2] <= 1'b0; cube[1][3][2] <= 1'b0; cube[2][3][2] <= 1'b0; cube[3][3][2] <= 1'b0; cube[4][3][2] <= 1'b0; cube[5][3][2] <= 1'b0; cube[6][3][2] <= 1'b0; cube[7][3][2] <= 1'b0; 
            cube[0][4][2] <= 1'b0; cube[1][4][2] <= 1'b0; cube[2][4][2] <= 1'b0; cube[3][4][2] <= 1'b0; cube[4][4][2] <= 1'b0; cube[5][4][2] <= 1'b0; cube[6][4][2] <= 1'b0; cube[7][4][2] <= 1'b0; 
            cube[0][5][2] <= 1'b0; cube[1][5][2] <= 1'b0; cube[2][5][2] <= 1'b0; cube[3][5][2] <= 1'b0; cube[4][5][2] <= 1'b0; cube[5][5][2] <= 1'b0; cube[6][5][2] <= 1'b0; cube[7][5][2] <= 1'b0; 
            cube[0][6][2] <= 1'b0; cube[1][6][2] <= 1'b0; cube[2][6][2] <= 1'b0; cube[3][6][2] <= 1'b0; cube[4][6][2] <= 1'b0; cube[5][6][2] <= 1'b0; cube[6][6][2] <= 1'b0; cube[7][6][2] <= 1'b0;
            cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
            cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0;
            cube[0][1][3] <= 1'b0; cube[1][1][3] <= 1'b0; cube[2][1][3] <= 1'b0; cube[3][1][3] <= 1'b0; cube[4][1][3] <= 1'b0; cube[5][1][3] <= 1'b0; cube[6][1][3] <= 1'b0; cube[7][1][3] <= 1'b0; 
            cube[0][2][3] <= 1'b0; cube[1][2][3] <= 1'b0; cube[2][2][3] <= 1'b0; cube[3][2][3] <= 1'b0; cube[4][2][3] <= 1'b0; cube[5][2][3] <= 1'b0; cube[6][2][3] <= 1'b0; cube[7][2][3] <= 1'b0; 
            cube[0][3][3] <= 1'b0; cube[1][3][3] <= 1'b0; cube[2][3][3] <= 1'b0; cube[3][3][3] <= 1'b0; cube[4][3][3] <= 1'b0; cube[5][3][3] <= 1'b0; cube[6][3][3] <= 1'b0; cube[7][3][3] <= 1'b0; 
            cube[0][4][3] <= 1'b0; cube[1][4][3] <= 1'b0; cube[2][4][3] <= 1'b0; cube[3][4][3] <= 1'b0; cube[4][4][3] <= 1'b0; cube[5][4][3] <= 1'b0; cube[6][4][3] <= 1'b0; cube[7][4][3] <= 1'b0; 
            cube[0][5][3] <= 1'b0; cube[1][5][3] <= 1'b0; cube[2][5][3] <= 1'b0; cube[3][5][3] <= 1'b0; cube[4][5][3] <= 1'b0; cube[5][5][3] <= 1'b0; cube[6][5][3] <= 1'b0; cube[7][5][3] <= 1'b0; 
            cube[0][6][3] <= 1'b0; cube[1][6][3] <= 1'b0; cube[2][6][3] <= 1'b0; cube[3][6][3] <= 1'b0; cube[4][6][3] <= 1'b0; cube[5][6][3] <= 1'b0; cube[6][6][3] <= 1'b0; cube[7][6][3] <= 1'b0;
            cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
            cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b0; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
            cube[0][1][4] <= 1'b0; cube[1][1][4] <= 1'b0; cube[2][1][4] <= 1'b0; cube[3][1][4] <= 1'b0; cube[4][1][4] <= 1'b0; cube[5][1][4] <= 1'b0; cube[6][1][4] <= 1'b0; cube[7][1][4] <= 1'b0; 
            cube[0][2][4] <= 1'b0; cube[1][2][4] <= 1'b0; cube[2][2][4] <= 1'b0; cube[3][2][4] <= 1'b0; cube[4][2][4] <= 1'b0; cube[5][2][4] <= 1'b0; cube[6][2][4] <= 1'b0; cube[7][2][4] <= 1'b0;
            cube[0][3][4] <= 1'b0; cube[1][3][4] <= 1'b0; cube[2][3][4] <= 1'b0; cube[3][3][4] <= 1'b0; cube[4][3][4] <= 1'b0; cube[5][3][4] <= 1'b0; cube[6][3][4] <= 1'b0; cube[7][3][4] <= 1'b0; 
            cube[0][4][4] <= 1'b0; cube[1][4][4] <= 1'b0; cube[2][4][4] <= 1'b0; cube[3][4][4] <= 1'b0; cube[4][4][4] <= 1'b0; cube[5][4][4] <= 1'b0; cube[6][4][4] <= 1'b0; cube[7][4][4] <= 1'b0; 
            cube[0][5][4] <= 1'b0; cube[1][5][4] <= 1'b0; cube[2][5][4] <= 1'b0; cube[3][5][4] <= 1'b0; cube[4][5][4] <= 1'b0; cube[5][5][4] <= 1'b0; cube[6][5][4] <= 1'b0; cube[7][5][4] <= 1'b0; 
            cube[0][6][4] <= 1'b0; cube[1][6][4] <= 1'b0; cube[2][6][4] <= 1'b0; cube[3][6][4] <= 1'b0; cube[4][6][4] <= 1'b0; cube[5][6][4] <= 1'b0; cube[6][6][4] <= 1'b0; cube[7][6][4] <= 1'b0; 
            cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b0; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
            cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0; 
            cube[0][1][5] <= 1'b0; cube[1][1][5] <= 1'b0; cube[2][1][5] <= 1'b0; cube[3][1][5] <= 1'b0; cube[4][1][5] <= 1'b0; cube[5][1][5] <= 1'b0; cube[6][1][5] <= 1'b0; cube[7][1][5] <= 1'b0;
            cube[0][2][5] <= 1'b0; cube[1][2][5] <= 1'b0; cube[2][2][5] <= 1'b0; cube[3][2][5] <= 1'b0; cube[4][2][5] <= 1'b0; cube[5][2][5] <= 1'b0; cube[6][2][5] <= 1'b0; cube[7][2][5] <= 1'b0; 
            cube[0][3][5] <= 1'b0; cube[1][3][5] <= 1'b0; cube[2][3][5] <= 1'b0; cube[3][3][5] <= 1'b0; cube[4][3][5] <= 1'b0; cube[5][3][5] <= 1'b0; cube[6][3][5] <= 1'b0; cube[7][3][5] <= 1'b0; 
            cube[0][4][5] <= 1'b0; cube[1][4][5] <= 1'b0; cube[2][4][5] <= 1'b0; cube[3][4][5] <= 1'b0; cube[4][4][5] <= 1'b0; cube[5][4][5] <= 1'b0; cube[6][4][5] <= 1'b0; cube[7][4][5] <= 1'b0; 
            cube[0][5][5] <= 1'b0; cube[1][5][5] <= 1'b0; cube[2][5][5] <= 1'b0; cube[3][5][5] <= 1'b0; cube[4][5][5] <= 1'b0; cube[5][5][5] <= 1'b0; cube[6][5][5] <= 1'b0; cube[7][5][5] <= 1'b0; 
            cube[0][6][5] <= 1'b0; cube[1][6][5] <= 1'b0; cube[2][6][5] <= 1'b0; cube[3][6][5] <= 1'b0; cube[4][6][5] <= 1'b0; cube[5][6][5] <= 1'b0; cube[6][6][5] <= 1'b0; cube[7][6][5] <= 1'b0; 
            cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
            cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0; 
            cube[0][1][6] <= 1'b0; cube[1][1][6] <= 1'b0; cube[2][1][6] <= 1'b0; cube[3][1][6] <= 1'b0; cube[4][1][6] <= 1'b0; cube[5][1][6] <= 1'b0; cube[6][1][6] <= 1'b0; cube[7][1][6] <= 1'b0; 
            cube[0][2][6] <= 1'b0; cube[1][2][6] <= 1'b0; cube[2][2][6] <= 1'b0; cube[3][2][6] <= 1'b0; cube[4][2][6] <= 1'b0; cube[5][2][6] <= 1'b0; cube[6][2][6] <= 1'b0; cube[7][2][6] <= 1'b0;
            cube[0][3][6] <= 1'b0; cube[1][3][6] <= 1'b0; cube[2][3][6] <= 1'b0; cube[3][3][6] <= 1'b0; cube[4][3][6] <= 1'b0; cube[5][3][6] <= 1'b0; cube[6][3][6] <= 1'b0; cube[7][3][6] <= 1'b0; 
            cube[0][4][6] <= 1'b0; cube[1][4][6] <= 1'b0; cube[2][4][6] <= 1'b0; cube[3][4][6] <= 1'b0; cube[4][4][6] <= 1'b0; cube[5][4][6] <= 1'b0; cube[6][4][6] <= 1'b0; cube[7][4][6] <= 1'b0; 
            cube[0][5][6] <= 1'b0; cube[1][5][6] <= 1'b0; cube[2][5][6] <= 1'b0; cube[3][5][6] <= 1'b0; cube[4][5][6] <= 1'b0; cube[5][5][6] <= 1'b0; cube[6][5][6] <= 1'b0; cube[7][5][6] <= 1'b0; 
            cube[0][6][6] <= 1'b0; cube[1][6][6] <= 1'b0; cube[2][6][6] <= 1'b0; cube[3][6][6] <= 1'b0; cube[4][6][6] <= 1'b0; cube[5][6][6] <= 1'b0; cube[6][6][6] <= 1'b0; cube[7][6][6] <= 1'b0; 
            cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
            cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b0; cube[4][0][7] <= 1'b0; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
            cube[0][1][7] <= 1'b0; cube[1][1][7] <= 1'b0; cube[2][1][7] <= 1'b0; cube[3][1][7] <= 1'b0; cube[4][1][7] <= 1'b0; cube[5][1][7] <= 1'b0; cube[6][1][7] <= 1'b0; cube[7][1][7] <= 1'b0;
            cube[0][2][7] <= 1'b0; cube[1][2][7] <= 1'b0; cube[2][2][7] <= 1'b0; cube[3][2][7] <= 1'b0; cube[4][2][7] <= 1'b0; cube[5][2][7] <= 1'b0; cube[6][2][7] <= 1'b0; cube[7][2][7] <= 1'b0;
            cube[0][3][7] <= 1'b0; cube[1][3][7] <= 1'b0; cube[2][3][7] <= 1'b0; cube[3][3][7] <= 1'b0; cube[4][3][7] <= 1'b0; cube[5][3][7] <= 1'b0; cube[6][3][7] <= 1'b0; cube[7][3][7] <= 1'b0;
            cube[0][4][7] <= 1'b0; cube[1][4][7] <= 1'b0; cube[2][4][7] <= 1'b0; cube[3][4][7] <= 1'b0; cube[4][4][7] <= 1'b0; cube[5][4][7] <= 1'b0; cube[6][4][7] <= 1'b0; cube[7][4][7] <= 1'b0;
            cube[0][5][7] <= 1'b0; cube[1][5][7] <= 1'b0; cube[2][5][7] <= 1'b0; cube[3][5][7] <= 1'b0; cube[4][5][7] <= 1'b0; cube[5][5][7] <= 1'b0; cube[6][5][7] <= 1'b0; cube[7][5][7] <= 1'b0;
            cube[0][6][7] <= 1'b0; cube[1][6][7] <= 1'b0; cube[2][6][7] <= 1'b0; cube[3][6][7] <= 1'b0; cube[4][6][7] <= 1'b0; cube[5][6][7] <= 1'b0; cube[6][6][7] <= 1'b0; cube[7][6][7] <= 1'b0;
            cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b0; cube[4][7][7] <= 1'b0; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
		end else begin
            if (been_ready && key_down[last_change] == 1'b1)begin
                if (!Pause) begin
                    A_pos_x <= next_A_pos_x;
                    A_pos_z <= next_A_pos_z;
                    B_pos_x <= next_B_pos_x;
                    B_pos_z <= next_B_pos_z;
                end
                Pause <= Next_Pause;
            end

            if (state == Play) begin
                cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b0; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b0; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b0; cube[4][7][7] <= 1'b0; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;

                cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b0; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b0; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0; 
                cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b0; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0; 
                cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0; 
                cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b0; cube[4][0][7] <= 1'b0; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0; 

                cube[A_pos_x + 1][0][A_pos_z] <= 1;
                cube[A_pos_x + 1][0][A_pos_z + 1] <= 1;
                cube[A_pos_x + 1][0][A_pos_z - 1] <= 1;
                cube[A_pos_x - 1][0][A_pos_z] <= 1;
                cube[A_pos_x - 1][0][A_pos_z + 1] <= 1;
                cube[A_pos_x - 1][0][A_pos_z - 1] <= 1;
                cube[A_pos_x][0][A_pos_z] <= 1;
                cube[A_pos_x][0][A_pos_z + 1] <= 1;
                cube[A_pos_x][0][A_pos_z - 1] <= 1;

                cube[A_pos_x][0][A_pos_z + 2] <= 0;
                cube[A_pos_x][0][A_pos_z - 2] <= 0;
                cube[A_pos_x - 1][0][A_pos_z + 2] <= 0;
                cube[A_pos_x - 1][0][A_pos_z - 2] <= 0;
                cube[A_pos_x + 1][0][A_pos_z + 2] <= 0;
                cube[A_pos_x + 1][0][A_pos_z - 2] <= 0;
                cube[A_pos_x - 2][0][A_pos_z] <= 0;
                cube[A_pos_x - 2][0][A_pos_z - 1] <= 0;
                cube[A_pos_x - 2][0][A_pos_z + 1] <= 0;
                cube[A_pos_x + 2][0][A_pos_z] <= 0;
                cube[A_pos_x + 2][0][A_pos_z - 1] <= 0;
                cube[A_pos_x + 2][0][A_pos_z + 1] <= 0;

                cube[B_pos_x + 1][7][B_pos_z] <= 1;
                cube[B_pos_x + 1][7][B_pos_z + 1] <= 1;
                cube[B_pos_x + 1][7][B_pos_z - 1] <= 1;
                cube[B_pos_x - 1][7][B_pos_z] <= 1;
                cube[B_pos_x - 1][7][B_pos_z + 1] <= 1;
                cube[B_pos_x - 1][7][B_pos_z - 1] <= 1;
                cube[B_pos_x][7][B_pos_z] <= 1;
                cube[B_pos_x][7][B_pos_z + 1] <= 1;
                cube[B_pos_x][7][B_pos_z - 1] <= 1;

                cube[B_pos_x][7][B_pos_z + 2] <= 0;
                cube[B_pos_x][7][B_pos_z - 2] <= 0;
                cube[B_pos_x - 1][7][B_pos_z + 2] <= 0;
                cube[B_pos_x - 1][7][B_pos_z - 2] <= 0;
                cube[B_pos_x + 1][7][B_pos_z + 2] <= 0;
                cube[B_pos_x + 1][7][B_pos_z - 2] <= 0;
                cube[B_pos_x - 2][7][B_pos_z] <= 0;
                cube[B_pos_x - 2][7][B_pos_z - 1] <= 0;
                cube[B_pos_x - 2][7][B_pos_z + 1] <= 0;
                cube[B_pos_x + 2][7][B_pos_z] <= 0;
                cube[B_pos_x + 2][7][B_pos_z - 1] <= 0;
                cube[B_pos_x + 2][7][B_pos_z + 1] <= 0;

                if (ball_pos_y == 3'd7 || ball_pos_y == 3'd0) begin
                    cube[ball_pos_x][ball_pos_y][ball_pos_z] <= 0;
                end
                else begin
                    cube[ball_pos_x][ball_pos_y][ball_pos_z] <= 1;
                end

                cube[prev_ball_pos_x][prev_ball_pos_y][prev_ball_pos_z] <= 0;

            end
            else begin
                case (A_score)
                    4'd0: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b1; cube[4][0][0] <= 1'b1; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b0; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b1; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b1; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b0; cube[5][0][4] <= 1'b1; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b1; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b1; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b1; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd1: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b1; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b0; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b1; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b1; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b1; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b1; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b1; cube[6][0][7] <= 1'b1; cube[7][0][7] <= 1'b0;
                    end
                    4'd2: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b0; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b1; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b1; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b1; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b1; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b1; cube[6][0][7] <= 1'b1; cube[7][0][7] <= 1'b0;
                    end
                    4'd3: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b0; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b1; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b1; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b1; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b1; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b1; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b1; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b1; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd4: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b0; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b1; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b1; cube[3][0][5] <= 1'b1; cube[4][0][5] <= 1'b1; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b1; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b1; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b0; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd5: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b1; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b1; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b1; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b1; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b1; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b1; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b1; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd6: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b1; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b1; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b1; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b1; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b1; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b1; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b1; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd7: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b1; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b1; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b0; cube[3][0][4] <= 1'b1; cube[4][0][4] <= 1'b0; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b1; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b1; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b0; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd8: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b1; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b1; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b1; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b1; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b1; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b1; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b1; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd9: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b1; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b1; cube[2][0][2] <= 1'b0; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b1; cube[2][0][3] <= 1'b0; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b1; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b1; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b1; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b0; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b1; cube[2][0][6] <= 1'b0; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b1; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    4'd10: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b1; cube[3][0][0] <= 1'b0; cube[4][0][0] <= 1'b0; cube[5][0][0] <= 1'b1; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b1; cube[5][0][1] <= 1'b0; cube[6][0][1] <= 1'b1; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b1; cube[5][0][2] <= 1'b0; cube[6][0][2] <= 1'b1; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b1; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b1; cube[5][0][3] <= 1'b0; cube[6][0][3] <= 1'b1; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b1; cube[5][0][4] <= 1'b0; cube[6][0][4] <= 1'b1; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b1; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b1; cube[5][0][5] <= 1'b0; cube[6][0][5] <= 1'b1; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b1; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b1; cube[5][0][6] <= 1'b0; cube[6][0][6] <= 1'b1; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b1; cube[3][0][7] <= 1'b0; cube[4][0][7] <= 1'b0; cube[5][0][7] <= 1'b1; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                    default: begin
                        cube[0][0][0] <= 1'b0; cube[1][0][0] <= 1'b0; cube[2][0][0] <= 1'b0; cube[3][0][0] <= 1'b1; cube[4][0][0] <= 1'b1; cube[5][0][0] <= 1'b0; cube[6][0][0] <= 1'b0; cube[7][0][0] <= 1'b0; 
                        cube[0][0][1] <= 1'b0; cube[1][0][1] <= 1'b0; cube[2][0][1] <= 1'b1; cube[3][0][1] <= 1'b0; cube[4][0][1] <= 1'b0; cube[5][0][1] <= 1'b1; cube[6][0][1] <= 1'b0; cube[7][0][1] <= 1'b0;
                        cube[0][0][2] <= 1'b0; cube[1][0][2] <= 1'b0; cube[2][0][2] <= 1'b1; cube[3][0][2] <= 1'b0; cube[4][0][2] <= 1'b0; cube[5][0][2] <= 1'b1; cube[6][0][2] <= 1'b0; cube[7][0][2] <= 1'b0; 
                        cube[0][0][3] <= 1'b0; cube[1][0][3] <= 1'b0; cube[2][0][3] <= 1'b1; cube[3][0][3] <= 1'b0; cube[4][0][3] <= 1'b0; cube[5][0][3] <= 1'b1; cube[6][0][3] <= 1'b0; cube[7][0][3] <= 1'b0; 
                        cube[0][0][4] <= 1'b0; cube[1][0][4] <= 1'b0; cube[2][0][4] <= 1'b1; cube[3][0][4] <= 1'b0; cube[4][0][4] <= 1'b0; cube[5][0][4] <= 1'b1; cube[6][0][4] <= 1'b0; cube[7][0][4] <= 1'b0; 
                        cube[0][0][5] <= 1'b0; cube[1][0][5] <= 1'b0; cube[2][0][5] <= 1'b1; cube[3][0][5] <= 1'b0; cube[4][0][5] <= 1'b0; cube[5][0][5] <= 1'b1; cube[6][0][5] <= 1'b0; cube[7][0][5] <= 1'b0;
                        cube[0][0][6] <= 1'b0; cube[1][0][6] <= 1'b0; cube[2][0][6] <= 1'b1; cube[3][0][6] <= 1'b0; cube[4][0][6] <= 1'b0; cube[5][0][6] <= 1'b1; cube[6][0][6] <= 1'b0; cube[7][0][6] <= 1'b0;
                        cube[0][0][7] <= 1'b0; cube[1][0][7] <= 1'b0; cube[2][0][7] <= 1'b0; cube[3][0][7] <= 1'b1; cube[4][0][7] <= 1'b1; cube[5][0][7] <= 1'b0; cube[6][0][7] <= 1'b0; cube[7][0][7] <= 1'b0;
                    end
                endcase

                case (B_score)
                    4'd0: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b1; cube[4][7][0] <= 1'b1; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b0; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b1; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b1; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b0; cube[5][7][4] <= 1'b1; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b1; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b1; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b1; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd1: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b1; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b1; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b1; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b1; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b1; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b1; cube[6][7][7] <= 1'b1; cube[7][7][7] <= 1'b0;
                    end
                    4'd2: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b1; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b1; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b1; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b1; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b1; cube[6][7][7] <= 1'b1; cube[7][7][7] <= 1'b0;
                    end
                    4'd3: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b1; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b1; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b1; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b1; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b1; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b1; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b1; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd4: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b0; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b1; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b1; cube[3][7][5] <= 1'b1; cube[4][7][5] <= 1'b1; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b1; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b1; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b0; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd5: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b1; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b1; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b1; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b1; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b1; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b1; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b1; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd6: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b1; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b1; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b1; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b1; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b1; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b1; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b1; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd7: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b1; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b1; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b1; cube[4][7][4] <= 1'b0; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b1; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b1; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b0; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd8: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b1; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b1; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b1; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b1; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b1; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b1; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b1; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd9: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b1; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b1; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b1; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b1; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b1; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b1; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b1; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b1; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b1; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    4'd10: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b1; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b0; cube[4][7][0] <= 1'b0; cube[5][7][0] <= 1'b1; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b1; cube[2][7][1] <= 1'b0; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b1; cube[5][7][1] <= 1'b0; cube[6][7][1] <= 1'b1; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b1; cube[2][7][2] <= 1'b0; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b1; cube[5][7][2] <= 1'b0; cube[6][7][2] <= 1'b1; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b1; cube[2][7][3] <= 1'b0; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b1; cube[5][7][3] <= 1'b0; cube[6][7][3] <= 1'b1; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b1; cube[2][7][4] <= 1'b0; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b1; cube[5][7][4] <= 1'b0; cube[6][7][4] <= 1'b1; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b1; cube[2][7][5] <= 1'b0; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b1; cube[5][7][5] <= 1'b0; cube[6][7][5] <= 1'b1; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b1; cube[2][7][6] <= 1'b0; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b1; cube[5][7][6] <= 1'b0; cube[6][7][6] <= 1'b1; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b1; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b0; cube[4][7][7] <= 1'b0; cube[5][7][7] <= 1'b1; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                    default: begin
                        cube[0][7][0] <= 1'b0; cube[1][7][0] <= 1'b0; cube[2][7][0] <= 1'b0; cube[3][7][0] <= 1'b1; cube[4][7][0] <= 1'b1; cube[5][7][0] <= 1'b0; cube[6][7][0] <= 1'b0; cube[7][7][0] <= 1'b0; 
                        cube[0][7][1] <= 1'b0; cube[1][7][1] <= 1'b0; cube[2][7][1] <= 1'b1; cube[3][7][1] <= 1'b0; cube[4][7][1] <= 1'b0; cube[5][7][1] <= 1'b1; cube[6][7][1] <= 1'b0; cube[7][7][1] <= 1'b0;
                        cube[0][7][2] <= 1'b0; cube[1][7][2] <= 1'b0; cube[2][7][2] <= 1'b1; cube[3][7][2] <= 1'b0; cube[4][7][2] <= 1'b0; cube[5][7][2] <= 1'b1; cube[6][7][2] <= 1'b0; cube[7][7][2] <= 1'b0; 
                        cube[0][7][3] <= 1'b0; cube[1][7][3] <= 1'b0; cube[2][7][3] <= 1'b1; cube[3][7][3] <= 1'b0; cube[4][7][3] <= 1'b0; cube[5][7][3] <= 1'b1; cube[6][7][3] <= 1'b0; cube[7][7][3] <= 1'b0; 
                        cube[0][7][4] <= 1'b0; cube[1][7][4] <= 1'b0; cube[2][7][4] <= 1'b1; cube[3][7][4] <= 1'b0; cube[4][7][4] <= 1'b0; cube[5][7][4] <= 1'b1; cube[6][7][4] <= 1'b0; cube[7][7][4] <= 1'b0; 
                        cube[0][7][5] <= 1'b0; cube[1][7][5] <= 1'b0; cube[2][7][5] <= 1'b1; cube[3][7][5] <= 1'b0; cube[4][7][5] <= 1'b0; cube[5][7][5] <= 1'b1; cube[6][7][5] <= 1'b0; cube[7][7][5] <= 1'b0;
                        cube[0][7][6] <= 1'b0; cube[1][7][6] <= 1'b0; cube[2][7][6] <= 1'b1; cube[3][7][6] <= 1'b0; cube[4][7][6] <= 1'b0; cube[5][7][6] <= 1'b1; cube[6][7][6] <= 1'b0; cube[7][7][6] <= 1'b0;
                        cube[0][7][7] <= 1'b0; cube[1][7][7] <= 1'b0; cube[2][7][7] <= 1'b0; cube[3][7][7] <= 1'b1; cube[4][7][7] <= 1'b1; cube[5][7][7] <= 1'b0; cube[6][7][7] <= 1'b0; cube[7][7][7] <= 1'b0;
                    end
                endcase
            end

            layer1 <= {
                cube[0][0][0], cube[1][0][0], cube[2][0][0], cube[3][0][0], cube[4][0][0], cube[5][0][0], cube[6][0][0], cube[7][0][0], 
                cube[0][1][0], cube[1][1][0], cube[2][1][0], cube[3][1][0], cube[4][1][0], cube[5][1][0], cube[6][1][0], cube[7][1][0], 
                cube[0][2][0], cube[1][2][0], cube[2][2][0], cube[3][2][0], cube[4][2][0], cube[5][2][0], cube[6][2][0], cube[7][2][0], 
                cube[0][3][0], cube[1][3][0], cube[2][3][0], cube[3][3][0], cube[4][3][0], cube[5][3][0], cube[6][3][0], cube[7][3][0], 
                cube[0][4][0], cube[1][4][0], cube[2][4][0], cube[3][4][0], cube[4][4][0], cube[5][4][0], cube[6][4][0], cube[7][4][0], 
                cube[0][5][0], cube[1][5][0], cube[2][5][0], cube[3][5][0], cube[4][5][0], cube[5][5][0], cube[6][5][0], cube[7][5][0], 
                cube[0][6][0], cube[1][6][0], cube[2][6][0], cube[3][6][0], cube[4][6][0], cube[5][6][0], cube[6][6][0], cube[7][6][0], 
                cube[0][7][0], cube[1][7][0], cube[2][7][0], cube[3][7][0], cube[4][7][0], cube[5][7][0], cube[6][7][0], cube[7][7][0]
            };
            
            layer2 <= {
                cube[0][0][1], cube[1][0][1], cube[2][0][1], cube[3][0][1], cube[4][0][1], cube[5][0][1], cube[6][0][1], cube[7][0][1], 
                cube[0][1][1], cube[1][1][1], cube[2][1][1], cube[3][1][1], cube[4][1][1], cube[5][1][1], cube[6][1][1], cube[7][1][1],
                cube[0][2][1], cube[1][2][1], cube[2][2][1], cube[3][2][1], cube[4][2][1], cube[5][2][1], cube[6][2][1], cube[7][2][1], 
                cube[0][3][1], cube[1][3][1], cube[2][3][1], cube[3][3][1], cube[4][3][1], cube[5][3][1], cube[6][3][1], cube[7][3][1], 
                cube[0][4][1], cube[1][4][1], cube[2][4][1], cube[3][4][1], cube[4][4][1], cube[5][4][1], cube[6][4][1], cube[7][4][1],
                cube[0][5][1], cube[1][5][1], cube[2][5][1], cube[3][5][1], cube[4][5][1], cube[5][5][1], cube[6][5][1], cube[7][5][1], 
                cube[0][6][1], cube[1][6][1], cube[2][6][1], cube[3][6][1], cube[4][6][1], cube[5][6][1], cube[6][6][1], cube[7][6][1], 
                cube[0][7][1], cube[1][7][1], cube[2][7][1], cube[3][7][1], cube[4][7][1], cube[5][7][1], cube[6][7][1], cube[7][7][1]
            };

            layer3 <= {
                cube[0][0][2], cube[1][0][2], cube[2][0][2], cube[3][0][2], cube[4][0][2], cube[5][0][2], cube[6][0][2], cube[7][0][2], 
                cube[0][1][2], cube[1][1][2], cube[2][1][2], cube[3][1][2], cube[4][1][2], cube[5][1][2], cube[6][1][2], cube[7][1][2], 
                cube[0][2][2], cube[1][2][2], cube[2][2][2], cube[3][2][2], cube[4][2][2], cube[5][2][2], cube[6][2][2], cube[7][2][2], 
                cube[0][3][2], cube[1][3][2], cube[2][3][2], cube[3][3][2], cube[4][3][2], cube[5][3][2], cube[6][3][2], cube[7][3][2], 
                cube[0][4][2], cube[1][4][2], cube[2][4][2], cube[3][4][2], cube[4][4][2], cube[5][4][2], cube[6][4][2], cube[7][4][2], 
                cube[0][5][2], cube[1][5][2], cube[2][5][2], cube[3][5][2], cube[4][5][2], cube[5][5][2], cube[6][5][2], cube[7][5][2], 
                cube[0][6][2], cube[1][6][2], cube[2][6][2], cube[3][6][2], cube[4][6][2], cube[5][6][2], cube[6][6][2], cube[7][6][2], 
                cube[0][7][2], cube[1][7][2], cube[2][7][2], cube[3][7][2], cube[4][7][2], cube[5][7][2], cube[6][7][2], cube[7][7][2]
            };

            layer4 <= {
                cube[0][0][3], cube[1][0][3], cube[2][0][3], cube[3][0][3], cube[4][0][3], cube[5][0][3], cube[6][0][3], cube[7][0][3],
                cube[0][1][3], cube[1][1][3], cube[2][1][3], cube[3][1][3], cube[4][1][3], cube[5][1][3], cube[6][1][3], cube[7][1][3],
                cube[0][2][3], cube[1][2][3], cube[2][2][3], cube[3][2][3], cube[4][2][3], cube[5][2][3], cube[6][2][3], cube[7][2][3], 
                cube[0][3][3], cube[1][3][3], cube[2][3][3], cube[3][3][3], cube[4][3][3], cube[5][3][3], cube[6][3][3], cube[7][3][3], 
                cube[0][4][3], cube[1][4][3], cube[2][4][3], cube[3][4][3], cube[4][4][3], cube[5][4][3], cube[6][4][3], cube[7][4][3], 
                cube[0][5][3], cube[1][5][3], cube[2][5][3], cube[3][5][3], cube[4][5][3], cube[5][5][3], cube[6][5][3], cube[7][5][3],
                cube[0][6][3], cube[1][6][3], cube[2][6][3], cube[3][6][3], cube[4][6][3], cube[5][6][3], cube[6][6][3], cube[7][6][3], 
                cube[0][7][3], cube[1][7][3], cube[2][7][3], cube[3][7][3], cube[4][7][3], cube[5][7][3], cube[6][7][3], cube[7][7][3]
            };

            layer5 <= {
                cube[0][0][4], cube[1][0][4], cube[2][0][4], cube[3][0][4], cube[4][0][4], cube[5][0][4], cube[6][0][4], cube[7][0][4],
                cube[0][1][4], cube[1][1][4], cube[2][1][4], cube[3][1][4], cube[4][1][4], cube[5][1][4], cube[6][1][4], cube[7][1][4], 
                cube[0][2][4], cube[1][2][4], cube[2][2][4], cube[3][2][4], cube[4][2][4], cube[5][2][4], cube[6][2][4], cube[7][2][4], 
                cube[0][3][4], cube[1][3][4], cube[2][3][4], cube[3][3][4], cube[4][3][4], cube[5][3][4], cube[6][3][4], cube[7][3][4],
                cube[0][4][4], cube[1][4][4], cube[2][4][4], cube[3][4][4], cube[4][4][4], cube[5][4][4], cube[6][4][4], cube[7][4][4], 
                cube[0][5][4], cube[1][5][4], cube[2][5][4], cube[3][5][4], cube[4][5][4], cube[5][5][4], cube[6][5][4], cube[7][5][4], 
                cube[0][6][4], cube[1][6][4], cube[2][6][4], cube[3][6][4], cube[4][6][4], cube[5][6][4], cube[6][6][4], cube[7][6][4], 
                cube[0][7][4], cube[1][7][4], cube[2][7][4], cube[3][7][4], cube[4][7][4], cube[5][7][4], cube[6][7][4], cube[7][7][4]
            };

            layer6 <= {
                cube[0][0][5], cube[1][0][5], cube[2][0][5], cube[3][0][5], cube[4][0][5], cube[5][0][5], cube[6][0][5], cube[7][0][5],
                cube[0][1][5], cube[1][1][5], cube[2][1][5], cube[3][1][5], cube[4][1][5], cube[5][1][5], cube[6][1][5], cube[7][1][5], 
                cube[0][2][5], cube[1][2][5], cube[2][2][5], cube[3][2][5], cube[4][2][5], cube[5][2][5], cube[6][2][5], cube[7][2][5], 
                cube[0][3][5], cube[1][3][5], cube[2][3][5], cube[3][3][5], cube[4][3][5], cube[5][3][5], cube[6][3][5], cube[7][3][5], 
                cube[0][4][5], cube[1][4][5], cube[2][4][5], cube[3][4][5], cube[4][4][5], cube[5][4][5], cube[6][4][5], cube[7][4][5],
                cube[0][5][5], cube[1][5][5], cube[2][5][5], cube[3][5][5], cube[4][5][5], cube[5][5][5], cube[6][5][5], cube[7][5][5], 
                cube[0][6][5], cube[1][6][5], cube[2][6][5], cube[3][6][5], cube[4][6][5], cube[5][6][5], cube[6][6][5], cube[7][6][5], 
                cube[0][7][5], cube[1][7][5], cube[2][7][5], cube[3][7][5], cube[4][7][5], cube[5][7][5], cube[6][7][5], cube[7][7][5] 
            };

            layer7 <= {
                cube[0][0][6], cube[1][0][6], cube[2][0][6], cube[3][0][6], cube[4][0][6], cube[5][0][6], cube[6][0][6], cube[7][0][6],
                cube[0][1][6], cube[1][1][6], cube[2][1][6], cube[3][1][6], cube[4][1][6], cube[5][1][6], cube[6][1][6], cube[7][1][6], 
                cube[0][2][6], cube[1][2][6], cube[2][2][6], cube[3][2][6], cube[4][2][6], cube[5][2][6], cube[6][2][6], cube[7][2][6], 
                cube[0][3][6], cube[1][3][6], cube[2][3][6], cube[3][3][6], cube[4][3][6], cube[5][3][6], cube[6][3][6], cube[7][3][6], 
                cube[0][4][6], cube[1][4][6], cube[2][4][6], cube[3][4][6], cube[4][4][6], cube[5][4][6], cube[6][4][6], cube[7][4][6],
                cube[0][5][6], cube[1][5][6], cube[2][5][6], cube[3][5][6], cube[4][5][6], cube[5][5][6], cube[6][5][6], cube[7][5][6], 
                cube[0][6][6], cube[1][6][6], cube[2][6][6], cube[3][6][6], cube[4][6][6], cube[5][6][6], cube[6][6][6], cube[7][6][6], 
                cube[0][7][6], cube[1][7][6], cube[2][7][6], cube[3][7][6], cube[4][7][6], cube[5][7][6], cube[6][7][6], cube[7][7][6] 
            };

            layer8 <= {
                cube[0][0][7], cube[1][0][7], cube[2][0][7], cube[3][0][7], cube[4][0][7], cube[5][0][7], cube[6][0][7], cube[7][0][7],
                cube[0][1][7], cube[1][1][7], cube[2][1][7], cube[3][1][7], cube[4][1][7], cube[5][1][7], cube[6][1][7], cube[7][1][7],
                cube[0][2][7], cube[1][2][7], cube[2][2][7], cube[3][2][7], cube[4][2][7], cube[5][2][7], cube[6][2][7], cube[7][2][7],
                cube[0][3][7], cube[1][3][7], cube[2][3][7], cube[3][3][7], cube[4][3][7], cube[5][3][7], cube[6][3][7], cube[7][3][7],
                cube[0][4][7], cube[1][4][7], cube[2][4][7], cube[3][4][7], cube[4][4][7], cube[5][4][7], cube[6][4][7], cube[7][4][7],
                cube[0][5][7], cube[1][5][7], cube[2][5][7], cube[3][5][7], cube[4][5][7], cube[5][5][7], cube[6][5][7], cube[7][5][7],
                cube[0][6][7], cube[1][6][7], cube[2][6][7], cube[3][6][7], cube[4][6][7], cube[5][6][7], cube[6][6][7], cube[7][6][7],
                cube[0][7][7], cube[1][7][7], cube[2][7][7], cube[3][7][7], cube[4][7][7], cube[5][7][7], cube[6][7][7], cube[7][7][7]
            }; 
		end
	end

    always @(*) begin
        case (last_change)
            A_Up: begin
                if (A_pos_z > 1'b1)
                    next_A_pos_z = A_pos_z - 1;
                else
                    next_A_pos_z = A_pos_z;

                next_A_pos_x = A_pos_x;
            end
            A_Down: begin
                if (A_pos_z < 3'd6)
                    next_A_pos_z = A_pos_z + 1;
                else
                    next_A_pos_z = A_pos_z;

                next_A_pos_x = A_pos_x;
            end
            A_Left: begin
                if (A_pos_x > 1'b1)
                    next_A_pos_x = A_pos_x - 1;
                else
                    next_A_pos_x = A_pos_x;

                next_A_pos_z = A_pos_z;
            end
            A_Right: begin
                if (A_pos_x < 3'd6)
                    next_A_pos_x = A_pos_x + 1;
                else
                    next_A_pos_x = A_pos_x;

                next_A_pos_z = A_pos_z;
            end
            default: begin
                next_A_pos_x = A_pos_x;
                next_A_pos_z = A_pos_z;
            end
        endcase
    end

    always @(*) begin
        case (last_change)
            B_Up: begin
                if (B_pos_z > 1'b1)
                    next_B_pos_z = B_pos_z - 1;
                else
                    next_B_pos_z = B_pos_z;

                next_B_pos_x = B_pos_x;
            end
            B_Down: begin
                if (B_pos_z < 3'd6)
                    next_B_pos_z = B_pos_z + 1;
                else
                    next_B_pos_z = B_pos_z;

                next_B_pos_x = B_pos_x;
            end
            B_Left: begin
                if (B_pos_x > 1'b1)
                    next_B_pos_x = B_pos_x - 1;
                else
                    next_B_pos_x = B_pos_x;

                next_B_pos_z = B_pos_z;
            end
            B_Right: begin
                if (B_pos_x < 3'd6)
                    next_B_pos_x = B_pos_x + 1;
                else
                    next_B_pos_x = B_pos_x;

                next_B_pos_z = B_pos_z;
            end
            default: begin
                next_B_pos_x = B_pos_x;
                next_B_pos_z = B_pos_z;
            end
        endcase
    end

    reg [2:0] abs_temp_x, abs_temp_z;

    always @(*) begin
        case (state)
            Play: begin
                if (ball_pos_y == 3'd0) begin // reach A
                    abs_temp_x = (ball_pos_x >= A_pos_x)? ball_pos_x - A_pos_x : A_pos_x - ball_pos_x;
                    abs_temp_z = (ball_pos_z >= A_pos_z)? ball_pos_z - A_pos_z : A_pos_z - ball_pos_z;
                    if (abs_temp_x > 1'b1 || abs_temp_z > 1'b1) begin // A dead
                        next_A_score = A_score;
                        next_B_score = B_score + 1'b1;
                        next_delta_x = 0;
                        next_delta_y = neg;
                        next_delta_z = 0;
                        next_ball_pos_x = 3'd4;
                        next_ball_pos_y = 3'd6;
                        next_ball_pos_z = 3'd4;
                        Next_state = ShowScore_1;
                    end
                    else begin // A catch
                        next_A_score = A_score;
                        next_B_score = B_score;
                        next_delta_y = pos;
                        next_ball_pos_y = ball_pos_y + 1;
                        next_ball_pos_x = A_pos_x;
                        next_ball_pos_z = A_pos_z;
                        next_delta_x = A_pos_x - ball_pos_x;
                        next_delta_z = A_pos_z - ball_pos_z;
                        Next_state = Play;
                    end

                end
                else if (ball_pos_y == 3'd7) begin // reach B
                    abs_temp_x = (ball_pos_x >= B_pos_x)? ball_pos_x - B_pos_x : B_pos_x - ball_pos_x;
                    abs_temp_z = (ball_pos_z >= B_pos_z)? ball_pos_z - B_pos_z : B_pos_z - ball_pos_z;
                    if ((abs_temp_x > 1'b1 || abs_temp_z > 1'b1)) begin // B dead
                        next_A_score = A_score + 1'b1;
                        next_B_score = B_score;
                        next_delta_x = 0;
                        next_delta_y = pos;
                        next_delta_z = 0;
                        next_ball_pos_x = 3'd4;
                        next_ball_pos_y = 3'd1;
                        next_ball_pos_z = 3'd4;
                        Next_state = ShowScore_1;
                    end
                    else begin // B catch
                        next_A_score = A_score;
                        next_B_score = B_score;
                        next_delta_y = neg;
                        next_ball_pos_y = ball_pos_y - 1;
                        next_ball_pos_x = B_pos_x;
                        next_ball_pos_z = B_pos_z;
                        next_delta_x = B_pos_x - ball_pos_x;
                        next_delta_z = B_pos_z - ball_pos_z;
                        Next_state = Play;
                    end
                    
                end
                else begin // in miidle
                    if (ball_pos_x == 3'b0 || ball_pos_x == 3'd7) begin
                        if (ball_pos_z == 3'b0 || ball_pos_z == 3'd7) begin
                            next_A_score = A_score;
                            next_B_score = B_score;
                            next_delta_x = neg * delta_x;
                            next_delta_y = delta_y;
                            next_delta_z = neg * delta_z;
                            next_ball_pos_x = ball_pos_x - delta_x;
                            next_ball_pos_y = ball_pos_y + delta_y;
                            next_ball_pos_z = ball_pos_z - delta_z;
                            Next_state = Play;
                        end
                        else begin
                            next_A_score = A_score;
                            next_B_score = B_score;
                            next_delta_x = neg * delta_x;
                            next_delta_y = delta_y;
                            next_delta_z = delta_z;
                            next_ball_pos_x = ball_pos_x - delta_x;
                            next_ball_pos_y = ball_pos_y + delta_y;
                            next_ball_pos_z = ball_pos_z + delta_z;
                            Next_state = Play;
                        end
                    end
                    else if (ball_pos_z == 3'b0 || ball_pos_z == 3'd7) begin
                        next_A_score = A_score;
                        next_B_score = B_score;
                        next_delta_x = delta_x;
                        next_delta_y = delta_y;
                        next_delta_z = neg * delta_z;
                        next_ball_pos_x = ball_pos_x + delta_x;
                        next_ball_pos_y = ball_pos_y + delta_y;
                        next_ball_pos_z = ball_pos_z - delta_z;
                        Next_state = Play;
                    end
                    else begin
                        next_A_score = A_score;
                        next_B_score = B_score;
                        next_ball_pos_x = ball_pos_x + delta_x;
                        next_ball_pos_y = ball_pos_y + delta_y;
                        next_ball_pos_z = ball_pos_z + delta_z;
                        next_delta_x = delta_x;
                        next_delta_y = delta_y;
                        next_delta_z = delta_z;
                        Next_state = Play;
                    end
                end
            end
            ShowScore_1: begin
                Next_state = ShowScore_2;
            end
            ShowScore_2: begin
                Next_state = Play;
            end
            default: 
                Next_state = Play;
        endcase
    end

    always @(*) begin
        if (A_score == 11 || B_score == 11)
            Next_Pause = 1;
        else
            Next_Pause = (last_change == Space) ? ~Pause : Pause;
    end

endmodule