`timescale 1ns / 1ps
// --------------------------------------------------------------------
// --------------------------------------------------------------------
// Module:top
// 
// Author: george
// 
// Description: top module of led cube
// 
// 
// --------------------------------------------------------------------
// Code Revision History :
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.0     |2021/01/11   |Initial ver
// --------------------------------------------------------------------
///////////////////////////////sample code : onepulse
module cube_top (
    clk,
    center,
    sw0,
    sw1,
    sw2,
    sclk_out,
    rclk_out,
    sdio_out,
    PS2_DATA,
    PS2_CLK
	);

    inout wire PS2_DATA;    
    inout wire PS2_CLK;
    input clk;
    input center;
    input sw0;
    input sw1;
    input sw2;
    output  sclk_out;
    output  rclk_out;
    output  sdio_out;

    wire clk_19;                            //1/2^17 clk = 2^27/2^17 = 2^10 = 1024 hz ~= 1ms   //digit period 
    clockDivider #(.n(19)) c19(clk, clk_19);//get 1/2^19 clk = 2^27/2^19 = 2^8 = 256 hz ~= 4ms //refresh period = digit period * 4

    wire debounced_center,onepulsed_center;
    debounce db(
        .pb(center),
        .clk(clk_19),
        .pb_debounce(debounced_center)
    );

    OnePulse op(
        .signal_single_pulse(onepulsed_center),
        .signal(debounced_center),
        .clock(clk_19)
    );

    reg [64-1:0] layer_1;
    reg [64-1:0] layer_2;
    reg [64-1:0] layer_3;
    reg [64-1:0] layer_4;
    reg [64-1:0] layer_5;
    reg [64-1:0] layer_6;
    reg [64-1:0] layer_7;
    reg [64-1:0] layer_8;

    wire [64-1:0] L1;
    wire [64-1:0] L2;
    wire [64-1:0] L3;
    wire [64-1:0] L4;
    wire [64-1:0] L5;
    wire [64-1:0] L6;
    wire [64-1:0] L7;
    wire [64-1:0] L8;
    
    Pong p(
        .clk(clk),
        .rst(debounced_center),
        .PS2_DATA(PS2_DATA),
        .PS2_CLK(PS2_CLK),
        .layer1(L1),
        .layer2(L2),
        .layer3(L3),
        .layer4(L4),
        .layer5(L5),
        .layer6(L6),
        .layer7(L7),
        .layer8(L8)
    );

   always@(*) begin
       if(sw0==1'b1) begin
           layer_1 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_00000000_00000000;
           layer_2 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_3 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_4 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_5 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_6 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_7 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           layer_8 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
       end
       else begin
           if(sw1==1'b1) begin
                layer_1 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
                layer_2 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_3 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_4 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_5 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_6 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_7 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                layer_8 = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;
           end
           else begin
               if(sw2==1'b1) begin
                    layer_1 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
                    layer_2 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_3 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_4 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_5 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_6 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_7 = 64'b10000001_00000000_00000000_00000000_00000000_00000000_00000000_10000001;
                    layer_8 = 64'b11111111_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
               end
               else begin
                    layer_1 = L1;
                    layer_2 = L2;
                    layer_3 = L3;
                    layer_4 = L4;
                    layer_5 = L5;
                    layer_6 = L6;
                    layer_7 = L7;
                    layer_8 = L8;
               end
           end
       end
   end 




    cube_scan cs
    (
        .clk_in(clk),			//系統clock
        .rst_n_in(onepulsed_center),		//系统reset，低位有效
        .layer_1(layer_1),	//單層LED第1排要顯示的數據
        .layer_2(layer_2),	//單層LED第2排要顯示的數據
        .layer_3(layer_3),	//單層LED第3排要顯示的數據
        .layer_4(layer_4),	//單層LED第4排要顯示的數據
        .layer_5(layer_5),	//單層LED第5排要顯示的數據
        .layer_6(layer_6),	//單層LED第6排要顯示的數據
        .layer_7(layer_7),	//單層LED第7排要顯示的數據
        .layer_8(layer_8),	//單層LED第8排要顯示的數據

        .sclk_out(sclk_out),		//74HC595的SCK腳位 //活塞 (SHCP) (SH)     //SRCLK//J2
        .rclk_out(rclk_out),		//74HC595的RCK腳位 //大平台 (STCP) (ST)   //RCLK//L2
        .sdio_out(sdio_out)		//74HC595的SER腳位 //資料 (DS)            //SER //J1
    );

endmodule
////////////////////////////////////////////////